module register_8(
    in,
    out,
    clk,
    rst,
    load
);
    input [7 : 0] in;
    output reg [7 : 0] out;
    input clk, rst;
    input load;

    always @(posedge clk, posedge rst) begin
        if (rst)
            out <= 8'b0000_0000;
        else
            if (load)
                out <= in;
    end

endmodule