`include "input_mux.v"
`include "weight_mux.v"
`include "bias_mux.v"
`include "PE.v"
`include "register.v"
`include "ReLU.v"
`include "counter.v"

module datapath(
    in,
    input_sel,
    reg_sel,
    weight_sel,
    bias_sel,
    clk,
    rst,
    reg_load,
    addr_count,
    addr_count_en,
    accuracy,
    acc_count_en,
    eql,
    expected
);
    input [62 * 8 - 1 : 0] in; //input from data_mem.v
    input input_sel, reg_sel;
    input [1 : 0] weight_sel, bias_sel; //weight and bias selection from controller.v
    input [30 - 1 : 0] reg_load; //register load from controller.v
    input clk, rst;
    output [9 : 0] addr_count; // label_mem.v, data_mem.v, and controller.v required
    input addr_count_en; //input signal from controller.v
    output [9 : 0] accuracy; //What we are looking for in Neural Processor
    input acc_count_en; //input signal from controller.v
    output eql; //output signal to controller.v
    input [3 : 0] expected; //What we expected from the input

    wire [7 : 0] bias_output [0 : 10 - 1];

    assign bias_output[0] = 8'b10000011;
    assign bias_output[1] = 8'b10101110;
    assign bias_output[2] = 8'b00100011;
    assign bias_output[3] = 8'b00000010;
    assign bias_output[4] = 8'b00010101;
    assign bias_output[5] = 8'b00000011;
    assign bias_output[6] = 8'b10011111;
    assign bias_output[7] = 8'b11000110;
    assign bias_output[8] = 8'b01010110;
    assign bias_output[9] = 8'b00000111;

    wire [7 : 0] bias_hidden [0: 30 - 1];

    assign bias_hidden[0] = 8'b00110100;
    assign bias_hidden[1] = 8'b00110110;
    assign bias_hidden[2] = 8'b10010001;
    assign bias_hidden[3] = 8'b11001110;
    assign bias_hidden[4] = 8'b11110100;
    assign bias_hidden[5] = 8'b11000111;
    assign bias_hidden[6] = 8'b10011110;
    assign bias_hidden[7] = 8'b11111111;
    assign bias_hidden[8] = 8'b10111000;
    assign bias_hidden[9] = 8'b11001111;
    assign bias_hidden[10] = 8'b01000011;
    assign bias_hidden[11] = 8'b11001001;
    assign bias_hidden[12] = 8'b00010000;
    assign bias_hidden[13] = 8'b00111001;
    assign bias_hidden[14]= 8'b10110010;
    assign bias_hidden[15] = 8'b11101010;
    assign bias_hidden[16] = 8'b11010111;
    assign bias_hidden[17] = 8'b11111111;
    assign bias_hidden[18] = 8'b10011101;
    assign bias_hidden[19] = 8'b10100001;
    assign bias_hidden[20] = 8'b11101111;
    assign bias_hidden[21] = 8'b01010011;
    assign bias_hidden[22] = 8'b00100101;
    assign bias_hidden[23] = 8'b11011100;
    assign bias_hidden[24] = 8'b00101101;
    assign bias_hidden[25] = 8'b10110110;
    assign bias_hidden[26] = 8'b00001011;
    assign bias_hidden[27] = 8'b11111011;
    assign bias_hidden[28] = 8'b11111111;
    assign bias_hidden[29] = 8'b11111111;

    wire [62 * 8 - 1 : 0] weight_hidden [0 : 30 - 1];
    
    assign weight_hidden[0] = 496'b10010011_00100001_00100111_00001111_10110011_10101001_00001110_10010110_01000101_10111010_00011100_11010010_10100000_11010110_10011110_10001011_11011011_00000001_10010011_10001001_10010010_10010001_01010000_00000001_11011001_11010111_10100100_10001111_01011110_00101101_00100111_01001010_01011000_10001110_10100000_00011010_00010010_11010011_10001001_00010100_11000001_10110000_10100010_01001101_01010001_00100111_00011000_00001100_01100011_10101101_10101011_10101101_01000101_10000100_00000100_10000011_10010110_00001111_00110011_00101000_10010110_10110011;
    assign weight_hidden[1] = 496'b10110000_10000100_00000100_00001111_10100110_10010001_00000001_10010000_00001111_10011011_10100000_10010100_10001111_00000100_00001100_00011000_00000000_00010011_10011011_00011111_10000110_11111111_10100001_10000001_10110000_00011010_00000100_10101111_10110011_11000000_00001100_00010000_00001010_10110001_10101010_10110000_00000011_10001101_00100011_00011101_00100001_00100011_00000010_00110010_00100010_00100100_00001100_00101001_00001110_00000011_10000011_10010011_00001111_00011000_00000011_00011111_00000001_00000001_10010100_10010101_00010110_10101011;
    assign weight_hidden[2] = 496'b11111111_10011100_11101001_00001110_10000110_00111011_00000111_11100001_10111011_10100010_00001010_00111111_00001100_00100110_00000111_10000111_01011010_10001101_10001010_01001001_00110001_10010001_10101010_10111110_00011100_00100000_00000100_00001000_10001100_01001010_00111111_00010011_10110001_10000001_10101100_00101011_10110011_10101010_10001011_10001000_00110000_00101110_11101001_00000000_00010111_00100011_00110101_00010101_00100000_11100001_10011001_00010111_00011111_00100010_01001111_10000001_00010000_11010010_10001110_00111011_10001000_11000010;
    assign weight_hidden[3] = 496'b10100110_00101111_00101111_00111100_11000100_00001101_10011001_00100111_00111111_00000010_10010011_00000000_10100110_00011001_11001110_10101001_00110110_01011000_10010001_00001111_10101100_00101000_10100001_00011101_00110000_00000101_10000001_10010100_10100000_10100111_00010001_10110101_10110001_00001001_10011000_11000101_10010101_00011001_00101101_10000011_10001101_11000011_00000110_00101011_10110101_01001011_10110001_10110101_10001011_01000000_10111100_10001111_00110000_10110100_10101010_00001100_00100001_10000101_00000111_00011011_10100100_11010001;
    assign weight_hidden[4] = 496'b10100111_10111000_00100110_00010100_10001101_10100011_10100110_00010100_10011001_10101110_00110111_11111011_10010001_00000110_10110100_00000010_10010100_10011011_00011101_10000101_00010110_00110001_00010111_10100101_00000101_10011100_00001010_10010101_00110110_00011110_00000110_10100001_11111111_10001100_10101111_10011101_01101101_10010111_10001010_00111111_10000110_10010101_00011101_00000110_10101100_00010001_00000010_00000100_00110011_00010011_00001111_10011000_00000101_00110110_00010111_00001010_00010001_00011101_10001000_00001110_00001111_10011100;
    assign weight_hidden[5] = 496'b10101000_10100000_10011111_10110111_00000110_10011100_10011010_10000101_10000011_10000101_00001001_10000011_00000000_00010110_10010001_00011001_11001101_00001110_00010001_00010011_00000101_10001101_10011011_00000010_00001110_00011111_10010111_10011001_10010111_10011010_10011101_00010100_00001101_00100011_00110101_10011110_10011010_01001001_00010000_00011111_10001111_00100010_00010001_00011010_00000101_00110011_10001010_00001110_00010010_10101100_00001110_10100110_00010001_10000010_00101001_10101100_00110001_10101111_11010000_00000001_00001110_00101000;
    assign weight_hidden[6] = 496'b00001111_10001111_10011000_10000101_00000101_10010010_10000001_10010000_10011011_00010110_10100010_10010101_10001110_00001110_10101101_11001101_01010000_10100000_11111111_10000010_00000011_00000101_10000110_10001111_10010011_01100010_10011001_10001000_00001001_00010001_10011010_11010000_10100010_10000010_00001101_00110111_10010110_00010000_10000110_01001000_01101110_00100001_10000001_10001101_10001101_10001000_11000001_00101010_10100010_00000000_00001101_00111001_10000111_01101011_10001011_10101111_00010011_00010010_10011100_00000000_10100001_11000110;
    assign weight_hidden[7] = 496'b00010110_10011100_10001100_00011100_11000110_01001100_00101101_01001101_10100010_00001110_11001001_11001100_10001111_10000110_01001000_01000001_11111111_10000111_00001111_10011000_10001001_10101011_00000110_00100110_10110101_00111001_00111010_00101101_10000011_11000011_10000101_01100011_10100111_10000001_10100110_10001111_10000011_10010111_10110000_10100101_11100100_10100000_00010100_10010010_00011101_10101110_10010000_10011111_00011010_00100000_10101110_10001101_10000110_11100100_00011001_10000011_10101101_10011010_10111001_00010011_10011110_10001010;
    assign weight_hidden[8] = 496'b11011001_00011000_10101100_10011001_00011011_00101010_00000101_11010001_00110111_10010011_10010111_10111001_00001111_00011101_00111001_10101010_00001111_00001111_10000010_00001000_10010110_10110000_00001101_10101011_10001110_00000101_10010100_10010001_00000000_10001100_00100101_10001101_00100111_00101010_00010100_10001001_10001000_00100011_00001010_00010010_00111101_01101011_00100000_00110101_10000110_10001010_11001000_10110001_11000111_11001010_10100010_00010010_00001100_00010110_10100101_00000010_00000101_10100010_00010101_10001111_10010000_11010011;
    assign weight_hidden[9] = 496'b10110110_10101011_10010011_10011100_10011010_11111111_00001100_10001110_10000011_00010001_11000100_01001000_10010100_11101100_01101010_11101000_11111111_00110001_11110010_00010111_10010110_11111001_00011100_10001011_11110001_10111000_10101110_00011110_00100000_00010001_00010011_01111111_01100001_01111111_01000000_00100101_11001001_10110101_11111111_10000100_10110011_01111111_11111111_10111110_00000000_00000110_01111111_00011101_10111000_00000110_10100100_01000101_10011111_00101000_10000111_00011110_01011110_00100000_10001101_00000000_00101100_01000001;
    assign weight_hidden[10] = 496'b10010010_10011011_10100001_00010100_10111000_00010000_00011100_10010000_10000011_10000010_10101011_01011001_00000101_00000111_00001110_00011000_00110001_00010010_00000101_00010001_10000001_10010010_10101110_10011001_10001101_10001000_10010001_00001110_10111101_00000110_00001110_01001001_00110111_10010111_00001111_10100110_11001011_10001101_10010101_00000110_00011101_00101010_11101101_10100100_00101011_00111100_00100111_10000111_00010001_11001011_00110001_11000100_00010110_00000001_00011011_10001010_10110100_00111110_00001110_10110111_00011111_00000011;
    assign weight_hidden[11] = 496'b00011011_10011110_10001000_10001110_10010001_10010011_00010010_00001100_00000000_00001000_10000111_00100011_10000100_00011111_00000001_00011000_00010110_10011101_11000000_01000010_10000011_10010000_10010000_00010110_10010011_00100110_10000010_00001100_10010010_10001101_01000001_00011111_10100000_11011001_10010110_10100111_00100111_00000010_00001000_10101111_10110110_10101101_10010011_10000101_00100001_00011011_00100111_00101110_10000100_10000010_10000010_10001001_10100010_10000011_10011010_10001011_10100000_10011101_10111000_00001000_00010101_11000101;
    assign weight_hidden[12] = 496'b10010011_10011100_10010100_00000010_00000010_00111101_00101000_00111111_00011000_10000110_00011100_00010111_10111011_00010100_10001000_00110111_00101000_10010000_01010010_00101001_00101011_10111100_10101011_00000000_00001111_10011010_00011111_00100101_00001011_10010010_00100001_11010110_10010111_10010101_00000101_00111000_00010011_00000001_00110110_00011001_00011000_10001001_11000111_10010110_10111100_11011001_10010111_10011100_10100100_00010011_10101010_10011000_10101000_10101001_10100101_10000101_10101001_00010010_10000101_00100100_10000001_00010100;
    assign weight_hidden[13] = 496'b00011001_10001010_10000010_10011001_00001011_10000110_00001100_00011100_10001001_00011000_10001010_00000110_10101100_00100001_01000010_10011101_10110010_00000100_00000000_00110011_10100010_00100010_10101101_00010000_10000001_10011011_10001011_00001001_10001001_00011000_10001010_00000101_00001001_10100000_00001100_00010010_00000011_00011110_00010101_10001111_10100000_10111101_10100010_00001010_00000111_00010100_00100011_00100011_10001101_00000100_00001001_00010010_10100011_00000010_10010101_10011000_00000111_00000000_00010001_10100011_00011001_00100000;
    assign weight_hidden[14] = 496'b00100001_10100010_10000011_10001000_00000000_00000101_00001000_10000100_10111100_10000011_10011100_00110111_00101011_00011110_00001101_10111001_11011000_00001010_11001011_10001001_10010011_10100101_00111000_10001000_10110011_01100010_00001000_00010100_00011001_10001101_10001010_10010101_11110010_01010010_00000011_00010011_00100001_00100001_10100000_00101001_10000011_00110001_01011110_00011001_10101001_10101110_10011000_00011100_00000011_00000001_10001111_10000001_00100101_11011001_00001101_10011100_00010010_10001110_00010011_10000001_00100001_00010010;
    assign weight_hidden[15] = 496'b00110110_00011000_10001001_00100100_01100000_00110001_10001111_10010100_10101001_00011010_00100110_10100000_10000111_10100010_10111100_11010101_11111001_11011101_00110010_00010010_10001011_00010010_10100110_00000010_10101011_00011011_00000100_10100110_10001010_10000110_10001011_10010011_10000101_10000001_10101100_00110000_11011101_10100011_11001011_10101000_10010100_10101000_11001101_10101100_00101011_00101111_00110110_10000100_10001000_10100110_00001011_10100010_10011001_10011111_00000111_00010100_10111101_00001011_00011111_00011010_11111000_00101001;
    assign weight_hidden[16] = 496'b00011010_00000000_00100010_00101010_00001000_01100011_00011010_00011111_10011010_10001010_10001110_11000101_11010110_10011110_10011010_00010110_00100101_10011101_10110100_00100110_00000101_10000010_10100000_00010010_10110101_00000111_11000000_10111100_00000011_10110010_00000101_10010001_11000110_10000011_10110101_10010100_00011110_10011001_00001010_00110111_10001000_10010110_10011101_00001000_00101111_00000011_10010000_00000110_00010110_10000011_00001000_00000100_00110110_00100011_00010011_10010111_00000111_10000001_10001111_00100111_11101010_00001001;
    assign weight_hidden[17] = 496'b00000000_10000001_00000000_10011011_00001110_10110100_10011111_10110001_10001000_00010001_11011000_00000111_00001110_00010001_10010000_10100101_10010001_00000000_10101011_10011111_10011011_10000010_00011110_10000100_00001010_10001110_00000110_00011111_00010000_10010111_00001010_00001101_00110011_00001101_00000001_00010111_00001111_00101011_00000000_10000001_00000100_00001100_10111001_00111101_10101011_00001110_10000111_00010001_10010111_11011101_00100000_00011011_10001111_00011001_00100111_11100010_00000010_00010111_10000111_00100111_10111001_10010000;
    assign weight_hidden[18] = 496'b00010101_10000001_00001111_10001100_00101000_10100010_10100110_10010001_00010001_00110001_11010110_00010011_10000100_10111011_10001000_10001010_00010101_00100110_00001000_10001111_10001010_10101110_00011111_10101010_00111011_10110010_10100111_10001010_10011011_10010111_00111111_10001001_10010100_00001001_10001000_00010100_10000111_11011110_00010001_10011000_10000001_00001100_00101101_10011000_00001111_10101010_10111010_10001111_00010000_00000101_00100000_11001011_00110000_00011000_10100000_10010101_10011101_00111011_10011001_01001110_00101101_10011000;
    assign weight_hidden[19] = 496'b00111110_11010110_00010100_10001000_10011110_10010000_00110110_00110000_10110001_00011110_00001000_00101110_10001010_10101000_10011001_00000001_00001010_00101111_10110101_11000111_00010011_10010101_10000111_00100000_10110101_10000011_00000011_00001000_00001100_10010100_10100110_00111110_10111001_00111001_10011101_10100111_10100001_10001100_11001101_00011111_10000111_01101010_10101011_10100111_10100100_10000011_10000001_00011001_10010001_00101101_00001001_00100101_00011010_10010001_10000100_10011000_00110111_00010101_00000101_10000100_00011101_00101010;
    assign weight_hidden[20] = 496'b10001000_10000011_10001101_10011001_00001111_00010001_00000001_00000111_00001111_00001001_10100001_10110111_10011100_00001100_00000111_00000010_00001110_10011100_00101100_01000100_00100010_00000010_10010000_00000111_10010011_01001010_10000101_00011010_10000101_00000110_00000000_00100100_10001101_00011000_00001001_10010011_00000001_00001000_00000011_10100010_10011100_00100101_10001101_10011011_00011111_10011100_00001111_10010011_10011111_00000011_11010011_00000100_10000101_10100011_10010111_00100101_11000010_10011101_10011010_00110000_00011001_11110010;
    assign weight_hidden[21] = 496'b10010111_00011101_10100011_00001000_00010001_10000110_10001000_10001111_00101101_00100110_10010000_00010111_00110101_00000100_10010110_00000011_00110111_10101000_00111000_10111001_00010010_00000011_00011011_01001000_00101011_10001101_00100001_00100001_10011110_00011101_11011101_01010110_00110100_10010111_00011011_10001001_10100010_10000001_11000100_00010111_00011000_00101110_00100000_11001110_01100101_10010001_00010110_01001100_00011010_10011100_10010011_00000010_00000000_10010100_00001100_00101110_10111110_10110011_00010011_00111011_11000001_11011100;
    assign weight_hidden[22] = 496'b10011010_10010110_10000001_10011010_00011000_10000001_10001100_10010000_00000011_10011000_00111111_10000110_00000110_00001010_10001001_10010110_00001001_00000011_01000111_10001000_10000101_10010001_00001001_00010110_00110101_11000101_10001000_10001000_00000101_00010000_00011011_10000110_00101111_10000101_10101000_00001101_00011111_10000010_10001001_00001000_00100010_10110011_10100001_00000000_00000000_00001101_10000100_00000000_00000011_10001010_00000011_10001010_11001010_00001111_10000001_10001001_00010100_10000111_00010100_00100000_00001100_10011100;
    assign weight_hidden[23] = 496'b10100111_01000110_10101011_00001111_10100111_00001100_10011100_10100100_00101010_00000000_00001110_10100101_00001000_10001100_10001101_11000101_10010011_10000101_00011101_00010101_10000010_00001010_00100111_00000010_10011011_00100111_10001110_00010101_10101010_00100101_10110010_00100010_00001010_00111111_00011100_00000100_00000111_00011001_10101010_10111100_10101011_10110010_10100001_00001110_10010001_00100000_11011111_10101100_10100010_10101110_00000001_00100010_10000110_00111000_00101001_00011000_00000010_00011010_10001010_00111011_10011010_00001111;
    assign weight_hidden[24] = 496'b00001110_10100000_10011111_00111000_00001001_10000110_10111001_00100100_10000010_10001111_00001010_10100010_00101111_01111111_11010111_00111111_10100110_10010010_10011011_00000101_10101111_01000000_10010110_00100100_11001001_01110111_00000101_00100000_10000011_10011000_10010100_00000100_00101010_10011000_11001111_11001101_10110101_10101001_11101111_10011010_00001010_00100111_00100100_00100100_00110000_01111111_00010111_00000111_10011011_10011000_00001000_10011001_00000010_11010000_00110001_10001000_00010101_10110000_00001111_10011111_10001010_00100000;
    assign weight_hidden[25] = 496'b10000100_11011110_10010110_00100000_00011101_10001100_00000111_10010010_11000110_00101110_10010001_00100010_00001100_10101101_10101000_00000011_11000011_00100000_10011000_10001000_00000100_10100101_00001001_10100010_00010101_00000110_00100100_00010100_10010111_00000110_01010100_11000100_10110011_00111111_10001000_00110111_10101100_10011010_10001101_00010110_00001000_00110111_00011010_10010000_01000010_00100111_00100010_00011100_10110000_10110001_00011001_10110011_00010110_11011100_10010110_10010001_00000000_10001110_00101001_00011111_10100000_00110001;
    assign weight_hidden[26] = 496'b00001000_00010110_10011000_10010011_10010111_11001011_00000111_10011100_00111011_00000111_10100000_00110000_00100111_10011100_00001000_00001000_00100110_00010000_10101101_10101000_00001010_10000001_00011001_10001111_00011110_10100101_10000001_10100000_10011100_10001011_10001010_00010100_00000001_10001010_10000100_10111001_10111100_10110011_10011111_10000011_00011110_00110101_00100100_10110100_10010011_10101111_10000001_00011010_00011111_00011111_10000101_00001110_10001010_00101001_10011110_10000001_00000011_00001001_00101000_00001000_10001000_10010011;
    assign weight_hidden[27] = 496'b10010011_00011100_01000000_00000011_00001000_00110000_00010101_10010011_11001001_00110111_10010010_00011010_10110111_10111010_00011000_10000111_10010011_10011001_00000000_10110000_00100000_10010011_10100001_10111001_10011001_00000001_01100011_10000011_00000110_11010111_10011000_00000011_00000001_10110111_10001001_10001111_11101110_00011011_10001111_10101101_00010001_00010111_10001000_00111101_10111010_10100010_00101101_10000111_10000100_00001011_00111101_01000000_10000111_10011011_00110111_10100010_10001100_00011111_00000101_10000100_10010101_10001010;
    assign weight_hidden[28] = 496'b10000100_10001010_10000010_10000111_00001100_10011010_10011001_10001110_10011110_10010001_10100100_11000000_10001001_10010000_10000001_00000100_00000011_10100101_00011001_00000110_00001001_00000010_10001111_00000000_10000100_10001000_00010011_00010100_10000011_10000100_10010000_00000100_00001010_00010001_00011110_10000010_10010000_00011001_00010001_10001010_00000100_00010001_10001001_00001100_00000011_00000010_00000110_00000000_10001111_00000101_10001011_00000001_00010110_10001101_10001010_00010000_10010000_00010111_10011110_10101101_10001000_11000010;
    assign weight_hidden[29] = 496'b10100010_00011011_00001010_10010010_00000100_00001100_00001000_10010000_00110110_10011100_00000001_10101111_00110011_10001001_00011110_01001111_00111110_10011111_00000000_10010011_00001000_00000101_00011010_00011000_10110000_10100110_00000111_00001011_00101011_00001101_10000111_00001001_00101100_00100111_10010001_00100010_10010011_10001011_00000101_11001011_10010110_00001100_00001001_00000111_10101001_10100010_10110111_10010111_10100011_10100111_10011011_00010100_10011011_10001100_10011100_10001010_10010100_10011100_10011001_10110011_00000010_10001000;

    wire [30 * 8 - 1 : 0] weight_output [0 : 10 - 1];

    assign weight_output[0] = 240'b00001100_10111010_10001010_10001101_10001010_10010000_10010000_00010001_00000001_00101111_00011101_00001100_00011001_10001011_00011101_10100011_10010111_10011110_10000001_00001011_00000011_10100100_10100111_10001110_00010101_00010000_00001101_10010101_00110110_10011001;
    assign weight_output[1] = 240'b00110110_10100000_10000110_10001000_00000101_10001101_00000100_10000100_00011100_10100111_00010001_00100110_00001100_10101010_00011100_10001001_00111111_10100110_10101100_10010010_10000101_00000110_00101000_00001111_10011110_00011100_00001000_00001100_00011010_10000100;
    assign weight_output[2] = 240'b10001101_10101000_10011111_00010111_10100101_00101000_10011010_00011111_10011110_00100010_00100100_00011101_00000110_00110101_10010001_10100110_10001110_00001011_10101101_10110110_00000100_10000011_10000111_10100101_10110010_10011000_10100010_00011110_10010010_10011110;
    assign weight_output[3] = 240'b10111000_11011000_00000101_10001001_11001011_00001101_10101001_11001100_00000110_10100100_10101000_00001101_00000001_10101010_00011000_00111000_10100101_00100010_00000011_11001011_00011100_00000110_10000011_10000101_00010010_00001011_00000101_00011000_10000001_00001011;
    assign weight_output[4] = 240'b10001101_00000011_10011001_00010001_00000100_10011010_10111011_10010000_10010001_01011010_10100011_11001100_01111010_10101110_00001101_10000101_00000011_10101101_10011011_00010001_10001101_10010011_00001001_10010100_10011100_10000110_10000111_00000100_10001000_10000010;
    assign weight_output[5] = 240'b10111100_10010100_00000011_00100110_00110010_10100110_01010101_11100110_10000010_10101001_10010001_10011001_10101001_10000100_00001101_10111010_00010010_00001001_00110100_10011001_10010111_00111110_10000001_10011110_10111001_00101011_10011001_10000011_00001011_10000110;
    assign weight_output[6] = 240'b00100001_10001000_00000110_10010111_00000001_00000001_00010101_00001010_00010000_10011101_10000100_00001110_10110100_00000111_10001011_10010001_10000011_00001111_00110110_00100110_00001011_00100011_00001101_00001100_00110000_00001110_00010111_10010101_10110001_10010011;
    assign weight_output[7] = 240'b00010010_01110100_00101110_01010101_00100000_00001000_10000100_00101011_10011111_00000110_10101110_10011101_10110010_00000110_00001000_00010001_00001011_00001100_10000110_00010110_00000001_10010011_00010000_00011000_01000000_00010101_00000011_10011001_10000001_00000000;
    assign weight_output[8] = 240'b10010101_11111111_10000011_10101010_00111111_10000010_10011011_00000010_10101010_00011011_10111011_10010111_10001011_00000001_10111110_10110001_10110110_10100001_10100000_00000001_10001000_10110000_10011001_00100110_10100011_10110110_10010010_10011111_10100011_00011110;
    assign weight_output[9] = 240'b10101101_01111111_11101110_10101011_10101111_00001110_10011101_10111000_00010010_11111111_00001000_00001100_11110000_11010000_00001000_10000001_10011010_10010100_00010101_00001101_00000011_00100010_00010111_00001100_11011111_10001001_00001100_00001011_10001011_00000011;

    wire [30 * 8 - 1 : 0] reg_hidden; //concatenation of output of 30 registers

    wire [62 * 8 - 1 : 0] input_out_mux [0 : 10 - 1];
    genvar i;
    generate
        for (i = 0 ; i < 10 ; i = i + 1)
        begin
            input_mux input_mux(
                .input_sel(input_sel),
                .reg_sel(reg_sel),
                .in(in),
                .reg_hid(reg_hidden),
                .out(input_out_mux[i])
            );
        end
    endgenerate

    wire [62 * 8 - 1:0] weight_out_mux [0 : 10 - 1];
    generate
        for (i = 0 ; i < 10 ; i = i + 1)
        begin
            weight_mux weight_mux(
                .weight_hid_i(weight_hidden[i]),
                .weight_hid_i_10(weight_hidden[i + 10]),
                .weight_hid_i_20(weight_hidden[i + 20]),
                .weight_out_i(weight_output[i]),
                .out(weight_out_mux[i]),
                .sel(weight_sel)
            );
        end
    endgenerate

    wire [8 - 1 : 0] bias_output_mux [0 : 10 - 1];
    generate
        for (i = 0 ; i < 10 ; i = i + 1)
        begin
            bias_mux bias_mux(
                .bias_hid_i(bias_hidden[i]),
                .bias_hid_i_10(bias_hidden[i + 10]),
                .bias_hid_i_20(bias_hidden[i + 20]),
                .bias_out_i(bias_output[i]),
                .out(bias_output_mux[i]),
                .sel(bias_sel)
            );
        end
    endgenerate

    wire [8 - 1 : 0] PE_out [0 : 10 - 1];
    generate
        for (i = 0 ; i < 10 ; i = i + 1)
        begin
            PE PE( 
                .bias(bias_output_mux[i]),
                .weight(weight_out_mux[i]),
                .in(input_out_mux[i]),
                .out(PE_out[i])
            );

        end
    endgenerate 

    // Three registers for each hidden layer
    wire [8 - 1 : 0] reg_hidden_out [0 : 30 - 1];
    generate
        for (i = 0 ; i < 10 ; i = i + 1)
        begin
            register reg_hid_1(
                .in(PE_out[i]),
                .out(reg_hidden_out[i]),
                .clk(clk),
                .rst(rst),
                .load(reg_load[i])
            );

            register reg_hid_2(
                .in(PE_out[i]),
                .out(reg_hidden_out[i + 10]),
                .clk(clk),
                .rst(rst),
                .load(reg_load[i + 10])
            );

            register reg_hid_3(
                .in(PE_out[i]),
                .out(reg_hidden_out[i + 20]),
                .clk(clk),
                .rst(rst),
                .load(reg_load[i + 20])
            );
            
        end
    endgenerate 


    assign reg_hidden = {reg_hidden_out[29], reg_hidden_out[28], reg_hidden_out[27], reg_hidden_out[26], reg_hidden_out[25], reg_hidden_out[24], 
    reg_hidden_out[23], reg_hidden_out[22], reg_hidden_out[21], reg_hidden_out[20], reg_hidden_out[19], reg_hidden_out[18], reg_hidden_out[17], 
    reg_hidden_out[16], reg_hidden_out[15], reg_hidden_out[14], reg_hidden_out[13], reg_hidden_out[12], reg_hidden_out[11], reg_hidden_out[10], 
    reg_hidden_out[9], reg_hidden_out[8], reg_hidden_out[7], reg_hidden_out[6], reg_hidden_out[5], reg_hidden_out[4], 
    reg_hidden_out[3], reg_hidden_out[2], reg_hidden_out[1], reg_hidden_out[0]};


    wire [3 : 0] prediction;
    ReLU ReLU(
        .in( {PE_out[9], PE_out[8], PE_out[7], PE_out[6], PE_out[5], PE_out[4], PE_out[3], PE_out[2], PE_out[1], PE_out[0]} ),    
        .enable(reg_sel),
        .max_val(prediction) 
    );


    counter Addr_counter(
        .clk(clk),
        .rst(rst),
        .cnt(addr_count),
        .cnten(addr_count_en)
    );

    counter Acc_counter(
        .clk(clk),
        .rst(rst),
        .cnt(accuracy),
        .cnten(acc_count_en)
    );

    assign eql = (prediction == expected) ? 1'b1 : 1'b0; 
endmodule

