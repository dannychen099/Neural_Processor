module bias_hidden_mem(
    bias_hidden0, bias_hidden1, bias_hidden2, bias_hidden3, bias_hidden4, bias_hidden5, bias_hidden6, bias_hidden7, bias_hidden8, bias_hidden9, bias_hidden10, bias_hidden11, bias_hidden12, bias_hidden13, bias_hidden14, bias_hidden15,
    bias_hidden16, bias_hidden17, bias_hidden18, bias_hidden19, bias_hidden20, bias_hidden21, bias_hidden22, bias_hidden23, bias_hidden24, bias_hidden25, bias_hidden26, bias_hidden27, bias_hidden28, bias_hidden29;
);
    output [7 : 0] bias_hidden0, bias_hidden1, bias_hidden2, bias_hidden3, bias_hidden4, bias_hidden5, bias_hidden6, bias_hidden7, bias_hidden8, bias_hidden9, bias_hidden10, bias_hidden11, bias_hidden12, bias_hidden13, bias_hidden14, bias_hidden15, bias_hidden16, bias_hidden17, bias_hidden18, bias_hidden19, bias_hidden20, bias_hidden21, bias_hidden22, bias_hidden23, bias_hidden24, bias_hidden25, bias_hidden26, bias_hidden27, bias_hidden28, bias_hidden29;

    assign bias_hidden0 = 8'b00110100
    assign bias_hidden1 = 8'b00110110
    assign bias_hidden2 = 8'b10010001
    assign bias_hidden3 = 8'b11001110
    assign bias_hidden4 = 8'b11110100
    assign bias_hidden5 = 8'b11000111
    assign bias_hidden6 = 8'b10011110
    assign bias_hidden7 = 8'b11111111
    assign bias_hidden8 = 8'b10111000
    assign bias_hidden9 = 8'b11001111
    assign bias_hidden10 = 8'b01000011
    assign bias_hidden11 = 8'b11001001
    assign bias_hidden12 = 8'b00010000
    assign bias_hidden13 = 8'b00111001
    assign bias_hidden14 = 8'b10110010
    assign bias_hidden15 = 8'b11101010
    assign bias_hidden16 = 8'b11010111
    assign bias_hidden17 = 8'b11111111
    assign bias_hidden18 = 8'b10011101
    assign bias_hidden19 = 8'b10100001
    assign bias_hidden20 = 8'b11101111
    assign bias_hidden21 = 8'b01010011
    assign bias_hidden22 = 8'b00100101
    assign bias_hidden23 = 8'b11011100
    assign bias_hidden24 = 8'b00101101
    assign bias_hidden25 = 8'b10110110
    assign bias_hidden26 = 8'b00001011
    assign bias_hidden27 = 8'b11111011
    assign bias_hidden28 = 8'b11111111
    assign bias_hidden29 = 8'b11111111